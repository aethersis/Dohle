.SUBCKT MN32xx Out1 Out2 Vdd In Vgg CP1 CP2 GND
C9          GND CP2 2.8N 
C10         GND CP1 2.8N 
C6          3 CP1 1.3P 
XT10        4 CP1 3 GND NMOSFET_0
XT11        3 Vgg 6 GND NMOSFET_0
XT9         7 Vgg 4 GND NMOSFET_0
C5          7 CP2 1.3P 
XT8         8 CP2 7 GND NMOSFET_0
XT13        9 Vgg 10 GND NMOSFET_0
C7          9 CP2 1.3P 
C4          11 CP1 1.3P 
XT6         12 CP1 11 GND NMOSFET_0
XT12        6 CP2 9 GND NMOSFET_0
XT7         11 Vgg 8 GND NMOSFET_0
C8          13 CP1 1.3P 
XT14        10 CP1 13 GND NMOSFET_0
XT16        14 CP2 Vdd GND NMOSFET_0
XT15        13 Vgg 14 GND NMOSFET_0
XT5         16 Vgg 12 GND NMOSFET_0
C3          16 CP2 1.3P 
C2          17 CP1 1.3P 
XT2         18 CP1 17 GND NMOSFET_0
C1          18 GND 1.3P 
XT4         19 CP2 16 GND NMOSFET_0
XT3         17 Vgg 19 GND NMOSFET_0
XT1         In CP2 18 GND NMOSFET_0
XT17        Vdd 9 Out1 GND NMOSFET_0
XT18        Vdd 13 Out2 GND NMOSFET_0

.ENDS

* CD4000 NMOS & PMOS TRANSISTORS
* TRANSISTOR MODELS ARE FROM LTSPICE GROUP MEMBER KCIN_MELNICK 
* SEE MESSAGE NUMBER 16897, HTTP://TECH.GROUPS.YAHOO.COM/GROUP/LTSPICE/ 
* NMOSFET DRAIN GATE SOURCE BULK 
.SUBCKT NMOSFET_0  1 2 3 4 
M1 1 2 3 4 CD4007N 
.ENDS 
* PMOSFET DRAIN GATE SOURCE BULK 
.SUBCKT PMOSFET 1 2 3 4 
M1 1 2 3 4 CD4007P 
.ENDS 
* 
.MODEL CD4007N NMOS ( 
+ LEVEL=1 VTO=1.44 KP=320U L=10U W=30U GAMMA=0 PHI=.6 LAMBDA=10M 
+ RD=23.2 RS=90.1 IS=16.64P CBD=2.0P CBS=2.0P CGSO=0.1P CGDO=0.1P 
+ PB=.8 TOX=1200N) 
* 
.MODEL CD4007P PMOS ( 
+ LEVEL=1 VTO=-1.2 KP=110U L=10U W=60U GAMMA=0 PHI=.6 LAMBDA=40M 
+ RD=21.2 RS=62.2 IS=16.64P CBD=4.0P CBS=4.0P CGSO=0.2P CGDO=0.2P 
+ PB=.8 TOX=1200N)


